.model m2n2222 npn is=19f bf=150 vaf=100 ikf=.18
+      ise=50p ne=2.5 br=7.5 var=6.4 ikr=12m
+      isc=8.7p nc=1.2 rb=50 re=0.4 rc=0.4 cje=26p
+      tf=0.5n cjc=11p tr=7n xtb=1.5 kf=0.032f af=1