.model m2n2907 pnp is=1.1p bf=200 nf=1.2 vaf=50
+      ikf=0.1 ise=13p ne=1.9 br=6 rc=0.6 cje=23p
+      vje=0.85 mje=1.25 tf=0.5n cjc=19p vjc=0.5
+      mjc=0.2 tr=34n xtb=1.5